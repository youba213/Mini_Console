----------------------------------------------------------------------------------
-- Company: UPMC
-- Engineer: Julien Denoulet
-- 
--	Package Casse-Briques
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package pong_pack is

	-- Definition d'un Type Tableau de Briques (2 Rangees de 9)
	type tableau is array (1 downto 0) of std_logic_vector(8 downto 0);


end pong_pack;
